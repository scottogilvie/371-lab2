library verilog;
use verilog.vl_types.all;
entity seg7Control_testbench is
end seg7Control_testbench;
