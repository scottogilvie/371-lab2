library verilog;
use verilog.vl_types.all;
entity fourFuncCalc_stated is
    generic(
        IDLE            : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        START_RUN       : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi1);
        START_STROBELO  : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi1, Hi0);
        START_STROBEHI  : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        START_DONE      : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi0, Hi0);
        COMPUTE_RUN     : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi0, Hi1);
        COMPUTE_LOAD1   : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi1, Hi0);
        COMPUTE_LOAD1_READ: vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi1, Hi1);
        COMPUTE_LOAD2   : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi0);
        COMPUTE_LOAD2_READ: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi1);
        COMPUTE_RESULT  : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi1, Hi0);
        COMPUTE_RESULT_LOAD: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi1, Hi1);
        COMPUTE_WRITE   : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi0, Hi0);
        COMPUTE_STROBELO: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi0, Hi1);
        COMPUTE_STROBEHI: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi0);
        COMPUTE_DONE    : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        DISPLAY         : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi0, Hi0);
        DISPLAY_READ    : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi0, Hi1);
        fnIdle          : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        fnStart         : vl_logic_vector(0 to 1) := (Hi0, Hi1);
        fnCompute       : vl_logic_vector(0 to 1) := (Hi1, Hi0);
        fnDisplay       : vl_logic_vector(0 to 1) := (Hi1, Hi1);
        opAdd           : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        opSub           : vl_logic_vector(0 to 1) := (Hi0, Hi1);
        opMul           : vl_logic_vector(0 to 1) := (Hi1, Hi0);
        opDiv           : vl_logic_vector(0 to 1) := (Hi1, Hi1)
    );
    port(
        ledr            : out    vl_logic_vector(9 downto 0);
        hex0            : out    vl_logic_vector(6 downto 0);
        hex1            : out    vl_logic_vector(6 downto 0);
        hex2            : out    vl_logic_vector(6 downto 0);
        hex3            : out    vl_logic_vector(6 downto 0);
        hex4            : out    vl_logic_vector(6 downto 0);
        hex5            : out    vl_logic_vector(6 downto 0);
        clk             : in     vl_logic;
        sw              : in     vl_logic_vector(9 downto 0);
        key             : in     vl_logic_vector(3 downto 0);
        rst             : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of IDLE : constant is 1;
    attribute mti_svvh_generic_type of START_RUN : constant is 1;
    attribute mti_svvh_generic_type of START_STROBELO : constant is 1;
    attribute mti_svvh_generic_type of START_STROBEHI : constant is 1;
    attribute mti_svvh_generic_type of START_DONE : constant is 1;
    attribute mti_svvh_generic_type of COMPUTE_RUN : constant is 1;
    attribute mti_svvh_generic_type of COMPUTE_LOAD1 : constant is 1;
    attribute mti_svvh_generic_type of COMPUTE_LOAD1_READ : constant is 1;
    attribute mti_svvh_generic_type of COMPUTE_LOAD2 : constant is 1;
    attribute mti_svvh_generic_type of COMPUTE_LOAD2_READ : constant is 1;
    attribute mti_svvh_generic_type of COMPUTE_RESULT : constant is 1;
    attribute mti_svvh_generic_type of COMPUTE_RESULT_LOAD : constant is 1;
    attribute mti_svvh_generic_type of COMPUTE_WRITE : constant is 1;
    attribute mti_svvh_generic_type of COMPUTE_STROBELO : constant is 1;
    attribute mti_svvh_generic_type of COMPUTE_STROBEHI : constant is 1;
    attribute mti_svvh_generic_type of COMPUTE_DONE : constant is 1;
    attribute mti_svvh_generic_type of DISPLAY : constant is 1;
    attribute mti_svvh_generic_type of DISPLAY_READ : constant is 1;
    attribute mti_svvh_generic_type of fnIdle : constant is 1;
    attribute mti_svvh_generic_type of fnStart : constant is 1;
    attribute mti_svvh_generic_type of fnCompute : constant is 1;
    attribute mti_svvh_generic_type of fnDisplay : constant is 1;
    attribute mti_svvh_generic_type of opAdd : constant is 1;
    attribute mti_svvh_generic_type of opSub : constant is 1;
    attribute mti_svvh_generic_type of opMul : constant is 1;
    attribute mti_svvh_generic_type of opDiv : constant is 1;
end fourFuncCalc_stated;
